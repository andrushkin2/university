-- megafunction wizard: %PARALLEL_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: parallel_add 

-- ============================================================
-- File Name: parallel_add0.vhd
-- Megafunction Name(s):
-- 			parallel_add
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 222 10/21/2009 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY parallel_add0 IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END parallel_add0;


ARCHITECTURE SYN OF parallel_add0 IS

--	type ALTERA_MF_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire2	: ALTERA_MF_LOGIC_2D (2 DOWNTO 0, 15 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (15 DOWNTO 0);

BEGIN
	sub_wire4    <= data0x(15 DOWNTO 0);
	sub_wire3    <= data1x(15 DOWNTO 0);
	result    <= sub_wire0(15 DOWNTO 0);
	sub_wire1    <= data2x(15 DOWNTO 0);
	sub_wire2(2, 0)    <= sub_wire1(0);
	sub_wire2(2, 1)    <= sub_wire1(1);
	sub_wire2(2, 2)    <= sub_wire1(2);
	sub_wire2(2, 3)    <= sub_wire1(3);
	sub_wire2(2, 4)    <= sub_wire1(4);
	sub_wire2(2, 5)    <= sub_wire1(5);
	sub_wire2(2, 6)    <= sub_wire1(6);
	sub_wire2(2, 7)    <= sub_wire1(7);
	sub_wire2(2, 8)    <= sub_wire1(8);
	sub_wire2(2, 9)    <= sub_wire1(9);
	sub_wire2(2, 10)    <= sub_wire1(10);
	sub_wire2(2, 11)    <= sub_wire1(11);
	sub_wire2(2, 12)    <= sub_wire1(12);
	sub_wire2(2, 13)    <= sub_wire1(13);
	sub_wire2(2, 14)    <= sub_wire1(14);
	sub_wire2(2, 15)    <= sub_wire1(15);
	sub_wire2(1, 0)    <= sub_wire3(0);
	sub_wire2(1, 1)    <= sub_wire3(1);
	sub_wire2(1, 2)    <= sub_wire3(2);
	sub_wire2(1, 3)    <= sub_wire3(3);
	sub_wire2(1, 4)    <= sub_wire3(4);
	sub_wire2(1, 5)    <= sub_wire3(5);
	sub_wire2(1, 6)    <= sub_wire3(6);
	sub_wire2(1, 7)    <= sub_wire3(7);
	sub_wire2(1, 8)    <= sub_wire3(8);
	sub_wire2(1, 9)    <= sub_wire3(9);
	sub_wire2(1, 10)    <= sub_wire3(10);
	sub_wire2(1, 11)    <= sub_wire3(11);
	sub_wire2(1, 12)    <= sub_wire3(12);
	sub_wire2(1, 13)    <= sub_wire3(13);
	sub_wire2(1, 14)    <= sub_wire3(14);
	sub_wire2(1, 15)    <= sub_wire3(15);
	sub_wire2(0, 0)    <= sub_wire4(0);
	sub_wire2(0, 1)    <= sub_wire4(1);
	sub_wire2(0, 2)    <= sub_wire4(2);
	sub_wire2(0, 3)    <= sub_wire4(3);
	sub_wire2(0, 4)    <= sub_wire4(4);
	sub_wire2(0, 5)    <= sub_wire4(5);
	sub_wire2(0, 6)    <= sub_wire4(6);
	sub_wire2(0, 7)    <= sub_wire4(7);
	sub_wire2(0, 8)    <= sub_wire4(8);
	sub_wire2(0, 9)    <= sub_wire4(9);
	sub_wire2(0, 10)    <= sub_wire4(10);
	sub_wire2(0, 11)    <= sub_wire4(11);
	sub_wire2(0, 12)    <= sub_wire4(12);
	sub_wire2(0, 13)    <= sub_wire4(13);
	sub_wire2(0, 14)    <= sub_wire4(14);
	sub_wire2(0, 15)    <= sub_wire4(15);

	parallel_add_component : parallel_add
	GENERIC MAP (
		msw_subtract => "NO",
		pipeline => 0,
		representation => "UNSIGNED",
		result_alignment => "LSB",
		shift => 0,
		size => 3,
		width => 16,
		widthr => 16,
		lpm_type => "parallel_add"
	)
	PORT MAP (
		data => sub_wire2,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "FLEX10K"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
-- Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
-- Retrieval info: CONSTANT: SHIFT NUMERIC "0"
-- Retrieval info: CONSTANT: SIZE NUMERIC "3"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTHR NUMERIC "16"
-- Retrieval info: USED_PORT: data0x 0 0 16 0 INPUT NODEFVAL "data0x[15..0]"
-- Retrieval info: USED_PORT: data1x 0 0 16 0 INPUT NODEFVAL "data1x[15..0]"
-- Retrieval info: USED_PORT: data2x 0 0 16 0 INPUT NODEFVAL "data2x[15..0]"
-- Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT NODEFVAL "result[15..0]"
-- Retrieval info: CONNECT: @data 1 2 16 0 data2x 0 0 16 0
-- Retrieval info: CONNECT: @data 1 1 16 0 data1x 0 0 16 0
-- Retrieval info: CONNECT: @data 1 0 16 0 data0x 0 0 16 0
-- Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add0.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add0.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add0.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add0.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL parallel_add0_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
